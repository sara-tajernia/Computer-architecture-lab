----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    05:16:55 03/15/2021 
-- Design Name: 
-- Module Name:    MUX4X1_con - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity MUX4X1_con is
    Port ( input  : in  STD_LOGIC_VECTOR (3 downto 0);
           select1 : in  STD_LOGIC_VECTOR (1 downto 0);
           output : out  STD_LOGIC);
end MUX4X1_con;

architecture Behavioral of MUX4X1_con is

begin
 output<=input(0) when select1="00" else
			input(1) when select1="01" else
			input(2) when select1="10" else
			input(3);
		

end Behavioral;

